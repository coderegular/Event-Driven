#2 AND(e,a,c)
#2 NOT(d,c)
#4 AND(f,d,b)
#2 OR(g,e,f)